
`default_nettype none
module main(
	input 	[9:0] 	SW,
	output 	[9:0] 	LEDR,
	output	[7:0]		HEX0,
	output	[7:0]		HEX1,
	output	[7:0]		HEX2
);

	// Part I
	//******************

		
	//seg7_dec SEG0(SW[3], SW[2], SW[1], SW[0], HEX0[7:0]);
	//******************
	
	
	// Part II
	//******************
	
	
	wire w_z;
	wire [3:0] w_m;
	wire [3:0] w_a;
	
	//comparator (i_v3, i_v2, i_v1, i_v0, o_z)
	comparator comp0 (SW[3], SW[2], SW[1], SW[0], w_z);
	
	//circuit_A (i_v2, i_v1, i_v0, o_a0, o_a1, o_a2)
	circuit_A circA (SW[2], SW[1], SW[0], w_a[0], w_a[1], w_a[2]);
	
	// circuit_B (i_z, o_seg[7:0])
	circuit_B circB(w_z, HEX1);
	
	// mux_2_1_1bit (i_a, i_b, i_sel, o_m)
	mux_2_1_1bit mux3 (SW[3], 0, 			w_z, w_m[3]);
	mux_2_1_1bit mux2 (SW[2], w_a[2], w_z, w_m[2]);
	mux_2_1_1bit mux1 (SW[1], w_a[1], w_z, w_m[1]);
	mux_2_1_1bit mux0 (SW[0], w_a[0], w_z, w_m[0]);

	// seg7_dec (i_m3, i_m2, i_m1, i_m0, o_seg[7:0])
	seg7_dec seg0 (w_m[3], w_m[2], w_m[1], w_m[0], HEX0);

	
	// bin_to_dec b2d(SW[3], SW[2], SW[1], SW[0], HEX0, HEX1); // test part 2 as a module
	

	
	//******************
	
	// Part III
	//******************
	
	/*
	//FA fa0 (SW[0], SW[1], SW[2], LEDR[1], LEDR[0]);  // test FA first
	
	//adder_4bit ([3:0]i_a, [3:0]i_b, i_cin, o_cout, [3:0]o_s)
	adder_4bit ad0 (SW[3:0], SW[7:4], SW[8], LEDR[4], LEDR[3:0]);
	*/
	
	//******************
	
	// Part IV
	//******************
	
	/*
	wire [3:0] w_s;
	wire w_cout;
	
	// adder_4bit ([3:0]i_a, [3:0]i_b, i_cin, o_cout, [3:0]o_s)
	adder_4bit add0 (SW[3:0], SW[7:4], SW[8], w_cout, w_s);
	
	// bin_to_dec_v2 (i_v3, i_v2, i_v1, i_v0, i_cin, [7:0]o_seg0, [7:0]o_seg1)
	bin_to_dec_v2 bin2dec0 (w_s[3], w_s[2], w_s[1], w_s[0], w_cout, HEX0, HEX1);
	
	// checkBCD ([3:0]i_a, [3:0]i_b, o_error)
	checkBCD cb0 (SW[3:0], SW[7:0], LEDR[9]);
	*/
	
	//******************
	
	// Part V
	//******************
	
	// TODO
	
	//******************
	
	// Part VI
	//******************
	
	// TODO
	
	//******************
	
	// Part VII (Mandatory for Graduate Students)
	//******************
	
	// TODO
	
	//******************

endmodule
