

`default_nettype none

module FSM_MicroInstr #
(
	parameter N = 4
)
(
	input clk,
	input reset,
	input [N-1:0] IB_BUS,
	
	output reg LatchA,
	output reg EnableA,
	output reg LatchB,
	output reg EnableALU,
	output reg AddSub,
	output reg EnableIN,
	output reg EnableOut,
	output reg LoadInstr,
	output reg EnableInstr,
	input [N-1:0]	ToInstr,
	output reg EnableCount
);

	reg [2:0] state, next_state;

	// States
	localparam [2:0] IDLE = 3'd0, PHASE_1 = 3'd1, PHASE_2 = 3'd2, PHASE_3 = 3'd3, PHASE_4 = 3'd4;

	// 1. State Register (sequential)
	always @(posedge clk) begin
		if(reset)
			state <= IDLE;
		else
			state <= next_state;
	end
	
	// 2. Next-State Logic (combinational)
	always @(*) begin
		
		next_state = state; // default: hold state
	
		case(state)
		
			IDLE: 
				begin		
					// Move to FETCH
					next_state = PHASE_1;
				end
			
			// FETCH Instruction
			PHASE_1:
				begin
					// Move to DECODE
					next_state = PHASE_2;
				end
			
			// DECODE Instruction	
			PHASE_2:
				begin
					// Move to EXECUTE A
					next_state = PHASE_3;
				end
				
			// EXECUTE A Instruction
			PHASE_3:
				begin
					// Move to EXECUTE B
					next_state = PHASE_4;
				end
			
			// EXECUTE B Instruction	
			PHASE_4:
				begin
					// Move to FETCH
					next_state = PHASE_1;
				end
				
			default: ;// None
		
		endcase
	end
	
	// 3. Output Logic (combinational)
	
	always @(*) begin
	
		// default all signals are zero
		LoadInstr 	= 1'b0;
		EnableInstr = 1'b0;
		LatchB 		= 1'b0;
		LatchA 		= 1'b0;
		EnableALU 	= 1'b0;
		EnableCount = 1'b0;
		AddSub		= 1'b0;
		EnableIN		= 1'b0;
		EnableA		= 1'b0;
		EnableOut	= 1'b0;
	
		case(state)
		
			IDLE: 
				begin
					// Initialize things if needed
				end
			
			// FETCH Instruction
			PHASE_1:
				begin
					// same sequence for all asm instructions
					LoadInstr = 1'b1;
				end
			
			// DECODE Instruction	
			PHASE_2:
				begin
					// same sequence for all asm instructions
					EnableCount = 1'b1;
					EnableInstr = 1'b1;
				end
				
			// EXECUTE Instruction
			PHASE_3:
				begin
					
					case(ToInstr)
						
						4'b0000: // NOP
							begin
								// do nothing
							end
							
						4'b0001: // ADD
							begin
								LatchB 		= 1'b1;
								EnableInstr = 1'b1;
							end
							
						4'b0010: // SUB
							begin
								LatchB 		= 1'b1;
								EnableInstr = 1'b1;
							end
							
						4'b0011: // OUT
							begin
								EnableOut 	= 1'b1;
								EnableA 		= 1'b1;
							end	
						
						4'b0100: // IN
							begin
								LatchA 	= 1'b1;
								EnableIN = 1'b1;
							end
						
						4'b0101: // LDA
							begin
								LatchA 		= 1'b1;
								EnableInstr = 1'b1;
							end
						
					endcase
					
				end
			
			// EXECUTE Instruction	
			PHASE_4:
				begin
					
					case(ToInstr)
						
						4'b0000: // NOP
							begin
								// do nothing
							end
							
						4'b0001: // ADD
							begin
								LatchA 		= 1'b1;
								EnableALU 	= 1'b1;
							end
							
						4'b0010: // SUB
							begin
								LatchA 		= 1'b1;
								EnableALU 	= 1'b1;
								AddSub 		= 1'b1;
							end
							
						4'b0011: // OUT
							begin
								// do nothing
							end
							
						4'b0100: // IN
							begin
								// do nothing
							end
							
						4'b0101: // LDA
							begin
								// do nothing
							end
						
					endcase
					
				end
		
		endcase
	end

endmodule

`default_nettype wire

